module usb_sequencer
  (
   input  clk,
   input  reset_n,
   input  rxf_n,
   input  txe_n,
   output rd_n,
   output wr_n, 
   output nibble_write_enable,
   output chunk_write_enable
   );

endmodule // usb_sequencer

   
   

   
